package Common_pkg is

  type led_state is (State0, State1, State2, State3, State4);

end package;

package body Common_pkg is

end package body;
